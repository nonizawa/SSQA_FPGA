module xorshift #(parameter integer WIDTH = 20, parameter integer TYPE  = 0) (prn, enable, clock, reset);

    output [WIDTH-1:0] prn;
    reg [WIDTH-1:0] prn;
    input enable, clock, reset;

    parameter integer REGWIDTH = (WIDTH <= 64) ? 64 : ((WIDTH <= 128) ? 128 : ((WIDTH <= 1024) ? 1024 : ((WIDTH <= 4096) ? 4096 : -1)));

    parameter integer TAP0 = (WIDTH <= 64) ? 1 : ((WIDTH <= 128) ? 1 : ((WIDTH <= 1024) ? 1 : ((WIDTH <= 4096) ? 5 : -1)));

    parameter integer TAP1 = (WIDTH <= 64) ? 1 : ((WIDTH <= 128) ? 7 : ((WIDTH <= 1024) ? 13 : ((WIDTH <= 4096) ? 22 : -1)));

    parameter integer TAP2 = (WIDTH <= 64) ? 54 : ((WIDTH <= 128) ? 1 : ((WIDTH <= 1024) ? 7 : ((WIDTH <= 4096) ? 27 : -1)));

    parameter SEED = ((WIDTH <= 64) && (TYPE == 0)) ? 64'b1010001110001101010000101101001000010001000111001100001110000110 :
                    (((WIDTH <= 64) && (TYPE == 1)) ? 64'b0010100001111001111011000001011001110011101010101101001100110111 :
                    (((WIDTH <= 64) && (TYPE == 2)) ? 64'b1011000101111010011110000000010111011101100001000111000011101010 :
                    (((WIDTH <= 64) && (TYPE == 3)) ? 64'b0010101010110010010000110000001110110011110010001011001000110110 :
                   (((WIDTH <= 128) && (TYPE == 0)) ? 128'b00111001111010110001100110011011011011010011000111100100100011001011111011111010100101010000111111111101011101010100011100110000 :
                   (((WIDTH <= 128) && (TYPE == 1)) ? 128'b10000010011000001111000001011111001101000101111100010010111011100111100000000000010010111111100111110111100101101110100010101101 :
                   (((WIDTH <= 128) && (TYPE == 2)) ? 128'b01100110001111110101001111000000100011110001000011011000000110111000001101001011000110101110100100101011101110001011101011110010 :
                   (((WIDTH <= 128) && (TYPE == 3)) ? 128'b00110110100111011001011101100000110011111110110100111100011000000001000111010000110110001011011011011101111101111110110000000111 :
                  (((WIDTH <= 1024) && (TYPE == 0)) ? 1024'b1101001010110100001101110010110010111100100111011001010001111010000001110101100010010000100001101010110100111011101100001010110010010110111100111010110001010010101010101110100001001001011101100111000001111001001101100010000101110001100110101011010010111000110001101000110010110000001010001101111110111110110001001111010101111110001001100110110110010000000011101000111110101011111111101011010101101000001100011011011110000001010010010100011100001000100110001101101000100001010101000001100101001110010100101001101101011010010011001100101000010011010000001001101101000100001111000000010100111010111000100100110100001011100000000111111111101011111011011000010100101101111001010011010110010101001100111010001111010111100010110010100101011000011010110100111000000001101110010110000000011000010010110000011000101100111000101011000100010010011101001101001111111010000000111100111101011100000100101101101001100101000110000001100100001001110100001101011001100110000101110001100111111010101111010111001100000000010010000110010001001100 :
                  (((WIDTH <= 1024) && (TYPE == 1)) ? 1024'b0001010010010111000010011111001101010000100100110010101001000000011100110000110000011111100101001101000101110100111111001110110111010101110111101010110010011111100100000101001000011101100011101100011101010101011000010111101101111001000111110010001001000001011111000110110000111100110100001001010101111010111100001111101100011101101010111101101000000011000011110010111000000010100101010011001111111000101111101010000100101000111001001011100111010001011010010110100100110010110010100111110111111011010111010111100110000111111111101001011100001111001000101000100110111010110010101000001100100010110000111110011000101011110000110000011100010000011111100000101100011101101001110011010010111110111110000000101111110001111001011111011010110100101100110010101100111011000010110001110001101110101100110111101010110111011100010101110100100111011000010010011110110110000100010000100101001100101111100011111011010010110000010010000100010001110011011101000011001100010010101100100110100010101101010000100110110000010010100001011110010000 :
                  (((WIDTH <= 1024) && (TYPE == 2)) ? 1024'b1000100001001001111000101110111010110101101101110100000001001100001011100111001101000100100010001110010010100000111000100111001011000000010100101101010010111000001100000010001101000010100011000111110100011000010000001110101111000000010010011111100001100111101101100100001111000111110001101100101001101001001110001100000111111101000010101101000110110001000110101101000001000100100001100110111001000101101111011010111011101101000101101001010001100001001001111001000000011110100010001111000000100011010011100111010000011001001011001110101101000000111001101000011110001100010010001100111000111101110011011000001010001001010001011111010011000011110011010011000111010000110100000111111011110111100000100011110110101111111110001000111101011110110100001000110001010010100111010110101000100111000001100101101000001011101011001011011011001001000100000100010011001101011100000010101001011001001101001010011100011001001001001100101000000101001110100001000011001000100101011001011110101001011000011011001101000001010011000101000001110100 :
                  (((WIDTH <= 1024) && (TYPE == 3)) ? 1024'b1110111001111100000110011101011101000101010010110110110101000001010111001011010101101100010101110110100011000010111010101010101101000111011100001000111100000111111011000011001011100010000011100000010100110010100111101110101010101001010101101111011000101110111000011101000101011100001010110101010111011110101011001010010000110110000100001100110011101011010111011000100000110100101101110101000000101111100111010010100100100101110001000000111111100001011000100111011011101101000100000001101111010000101101010111101100100110011101110010001010110011111010000011101111101001111101110001011111000011100111110110110100110111001000100010111111001100101001001000110110010010111011101001100111000111010001111101001011100000000110000100100001111111000110010100011000010111001101011000100011011111110110011010101111010100100110111110110100011101111100000100010111011101100111110101010110100101011111111000000111001011011100001110010011100011000011011000011100000010011010111000101110001011011000011111101011111111111111111010001101001011 :
                  (((WIDTH <= 4096) && (TYPE == 0)) ? 4096'b1011011010110101100000100110001111111000111100001000010100110110100001001011110010000111011010101011010010111000000110000100000000110011010010110111010101001101000011100011011010000000011000010011000110010010101111101001100110101000111011100001010100001000100010101100100001011000101110100101110100001010011111110000001101100000010110001100101100001001001110101101010011111001111001001010100001110110110110110110010111010100011101101100111010011100000100100001001100110001010101010101011110001000011111100111001010000111110000001100111111101100111111101111010100010110011000001100101001110100000111001010111110011111100011110010110101000010001110101100010110101100111100111001001000110000001101010001010101100110000101010011001010111110011110111010011010100101111000010000100010110011110110011100100000011110111001010110000110111011111101111001101111010000101000000001111001001010101010011111100111101011000011000010111100010011111101101011010100010001010111001110100110110011010001010101110010111101011011100101100001101111011000111010101000101000110110011100111010000000010101001101111000101111110110100111011101101011101111100101000010010101001110000001001100011011001110010100100111100110011010000011001010011101010010001000010001010100111010110101111101000110110111010001011110100100011011100111101100100010000100110001100010101000110110100000100100001110011100011100101100000110110001010011110100001101000101100001111011011011001100001010111011001110011100100100100101011001111001110110110101011100100001000011010100100001011111010101100001111101000000000101110000001101010111000110000111000010101010101000101111101011000011001001011111110011011011001001100100100110001101110101111110100001010101111100101011101010111011000000001111001111001011000100101110100110110101110111011010101011100111100111111110000011001101001110000011010011100001100101101100000010001001111000011100010111011000111111111100011111101010100101110000101111001001101001000111110010011011110101010011011101100110101010111111101000100011011011100100101010100101011110000001010010010111110011110011010001101001101110100100011011000001110000100000000011000110100001110001001100100000000101001101001000100110100001001010100000101001110011001001100110000101000010000000100110101010111000001010000010000110100001010010100110100001000000111000001001100101011001011111000110010101001101101100011001100111110110100001000011111001100110000011110001101110011100100000110110010001100100000100101010011010011000001110000100011011101110100111110110111011000000011011010011010011110110011000110011101101101110111110100000010011111001110111011011101101101101001110111001111100110111010101001100111100000100101111001111010111001010110011000100100101110100000100101010110110111010100001001100001001101000011011011010101100110110010011010010011010011101110001100001100110000101100010101101101110000010001000011111111001101101111001101100000001101000100100000000111010100100100010010100010101100010010001001000100110111011111111011011100100100000111101010010001001101101101101000010011101101011010101100111010111001001011000010100100101101110110101111110001101001001110101000101010010010010011101100100001110100010100010100000101000001010000010000000100111111100011100100000100000010000100001010011110110111011101111010101111001000011000110110001001111100011100011100100001110101000000101011000000111100011011010010101101110100010001100001110101010100110001010011100010110101011010101000010100010011100110100100100011000110011100101100010111001011101111001100010010100101110011010100100011100001011110110001010101100011111110011111001110000101011001110000100111001001100000110111101101010000101010111100101000011011110101010111101101101101110000110001100100000010101010110010000000110111101110001110001000101001101111101001011110011011010111010100011001111101011001010101100010000010100101100111101010100100110110010100111001110100001101100100110000100100111010011111100000001011000000011011110101100010010010111001101110000010101001100111110000001010111001110000000011001110110011101001001101011110001011001111001110101100011011000011010 :
                  (((WIDTH <= 4096) && (TYPE == 1)) ? 4096'b1011111000100111101001010000101110011001001100101011000111000010111111000011000000000101011101001111010000011110100000001001111111111001011111011010111011110100110000111110110000011010100100101000111101010010100001110011110010111110110110011010111000010101001000100000111111011010000010001001000101100101111000001111011011100010110010111100111011110111110111110100100011111001010110100001100011100111110100000111100101001001110110011011101001111000111011100010011000111011111110100011000110010010001110010110110000011100001011000010101111100100100011101100111010101000110101001010101110100111010111111110100101000010111100001011001101100111101100001011001001111110111001110011110001110110001111101110011110111010001000100010000101010010100110011110010010110001000010101111110001111111110001001110010110010000111010011101010001001100010101000000111001000111001001110001101001001100111000001011010001100000100111111011101110001001011011100001110100011100100000001000001111111100001010000110101000001110011101010110100011110111100001011110011001100111101011010011000010100101010011110000110011101000001010101010011010100000100111110011011111001111100001011100010001011000100100000001000010000001001001000111010100011001111000100001111111110111010101000101010100011011101111101001111111111001011010110001010101111000000010001011001000011100000101000001001110011000100110000110101110000111111100011111111101100111000100110101011101010011010000001100110011000110101100111100011001110111010110010110001010000100100111001011011011101111010100001101011001100111000001101110001000000000100000000011100110110111011101011110110001111101101101010001101111101100110010000000011111111101101001111010110000000011000011111111000000010000000110110100011000011011101100000110000001001001011111101001010101011101111010101110111000000101111101001110111001101110010111001001100001110001100111100101110011110011101111001011100110010110011001101010010010100011011000001111001001101000101100010001011010100110000011110011011100001000010010010101010010100100000001101111111111101100110010100101110101011010100101011100100000001110000011011111100101000110111100001100001100101011100111011101011100010000111100011111000100100111011110111101000100011111110101100110000010011001100011110011011000101001010010011111110111111110000010101001000001101010110001100011111001010111010000100101100110001000101110000000001101001011111111110100010000111011001010000110101101100011100000011101001010000111010110011010000100101000110110101000010001101100010001010000101001011000010011001001011000111001000001001100111101010001101001010101001110110110011100110100010001000100000001001101100100001010110101101101110011100100101010101110000010101000100011000110110000011100000110000010001101110011111011110100001101101100011010001101010011101001011011100111111010101001101001011001101000000011101001001110111011110110010111010001101101111000110100100111111011101110010111100101110011111011100000110111000111101000101101101111101100000111010000000101000111101000010101110010111011001101010010101001111110010010101010101000001010100000101000001111100001001111000100011110011111110100011010011011110101100010010001101100001000001001001011101001010101110101000100100111111011001101110011000001010111000100011001101011011001001101101001010100111100111011001100000001100101011111110111011110000000110011110000011001111110000101011010000111010000101011000101001001101001000010010110111100110111101100100110010011111100101101101010111001110011100100001101110101111110010101010000110110110001010111000111100010111111010011010101000011011011100100001011001100000100001101001011100001111100000110011011110010111101001111010100011100110100001100000000011111101111000001100001100111000101100001111000110010101101011100100011001000101111111011000110011011110111101011010101011101001000000100001111100000011100000110010011010000100011101100011101100010010001110011101100001010000111001011100011011011000000100011010011010101111001010101110001110110101011110011111011111110010000101010001100000001001110100000011111000101000011101110000011000010001001110111 :
                  (((WIDTH <= 4096) && (TYPE == 2)) ? 4096'b1011000010100000101100000001001001101011011001000111100100011001000100011101110110001100011001101111101111101000100100101000010011000011010001100011010111110110111001111011110101001001111111101000110101101111110100011001101100110111001011000010000010100110111000011100001111111110101110110100010000100001101010000101000101110110100111001110010010000110111101011110000110010010011111110111010101000100011100100110101110110001011101101000011111101100001010110111001011010101101101110011100110000111010000010011010110110111100101001000111101110001111101101101100010101110000101100111111110011110100101110000110110010001111011100100101101011111110100111100000111011101010001011011110001110100110000000001010000110000110100101101011011010101100110001100010111011010001111111101110110111011101111111111111111001110100100000111001111010001011001101010111101001011110110011010000010111111100010010101011000010000110000001011001011000001001000101001001000100010010010001011101001100110100110000110010111000101001101100000000010101100000001101000010110011101010001010101001101000010101101101000001111010101111111010101001100111011000110111001111100101100001011110100001111000010111101111101010000101111010110111000111011111001100111100111111001100110110011000101101000101011111110011111100011111101100110111110000101110100101101001101000101001010001001001100101010001011011011010111110101100010001101101001000001110000011101100110001000001001001001101000001010111011000111111110000011001101101000110010110100101111001110100001111100111111101100110101100000011010100000010110010100100001011000100010000101110110010000110011011111011010101110010111011100111100100011111101011100101110011000011011100110000010011100111110011101011101100011011010011101110101100000011010000111011101011101100111110100001000011000111101110101011011001011010110111001101110010001101001110000110010001101110111011101111110111001110110111001100010011010100111000011101010111110110001110100110000011001011000000101010011101000001111100001101101101000011011110000101110001111110000101110000000100000011011110101000010001010111110000011111110110000000111000010111000100101011000101000100111010110101101100011001010110110011101111101000000111110001101110110000010001111101101100101100110000001011111011011010100100111000000000111010110101001110110101011110011010010010111101010001010010100011100001000101001001111101011100000010101110101111001101100001110000010000001100110100000101101010100011010110010110010001001101110001010110001101100011001110110110100000000010110100010111101110110010001010000001000010101010011001111001001110000110110011010111010110110111111000010010110100110101001000101011110100011001100010111101101000110101010100000010011111011000011011101011001010010010000010010001010101101011101101110001001010101011101000101010111010010111001001111100111010001001010111000011111100100010100110111100001010100100010111010100010011011111101100010111100001110010111011111011110011001110010010110101010100101110101110101110000111110001110010100101110111110111000110100011001011010000010011010000010001111000100110011000101111110100101110000000001110010101111110101001001011011000100011101001101000100101101010001110010001111010110010100111010000111000010001110111111110101101010110011010011010000011001000010101010101011010100011110001010111111101110101101101110110100110000101111111011011011010001001010001100011111111010111110000011001101000111110100010010011100010100011000000110001101110100010011110011101000110111111110101110000010110010001101100100011101100001000011000010100001101011101110000000110011011001100110001100110100000110010010011110110010100100001100110101011001010000011000100100011100101100011111010100001001110111001110000000010111001101110101111001111101001111100001010110110111100000011011000011100001010110001100000000111000010100001011100100111100011001011101100011110100000101110010000000000001101001110100001101000001000101101100111000011000001100101110011101000010011111111100101100101110101001111101101101111111111100110101101010100100100001101100110010110010100010001111101110101011001110111010 :
                  (((WIDTH <= 4096) && (TYPE == 3)) ? 4096'b1110110110100110001011001100011000100101011011111000101110100011010010100100001010111110011001011110001011111011011110010101101000101101111101101010111011000000011101111010010000011110001010001110011001010000101011000001011001001111110101001000100110001100101000000110101000110100000110100001110111011110000110101111000010110011001101011100011100011100100010110100000000011101100101001101000000011110000110101010010011111000000000000001000110011000111011010100100100001001110010101010111101001111100001011110100111010111110000000110110110010110001101100010000110010100110010010000111110100101011011001011011011001011010111111111011010010001101010000001110001100011100010101010111000000001010110100000000001100100010100110101001101100001001000100000001011100010001101110010110101000011110000001110110000100101010001110000101011011001000010001101100010101111000001101010011010100100110001101000100011100011001011100010001100010101001110100000110101110001001101101010110000111001011011001001011101110000100111110110101001001010001101110001111110100110101000110011000001111101011111101000100111000110011101110100101011001011110011101101101001011100010100100110011001010000110100011011011111111110110011010011010000111111100010010000110100100010011111100111000000010001100101000001100111010100000110000011111110001110010110101100011111001110001100101111000110110101101101101010100101111010011000000011000110000111000100001000001001001001000001010100100000100001100011110001000100111111010110011101110101111100000010000101011110100000100110011011101100000010101111011111010100011110110110001111110110001110101011111000101100010111011111000101001111110011100101011010111010100010001001111010111000001011001111101101010100000101001111110100101110010010101000001001100100001000000110110001100000111101000101111011100101100100100101100000001000100000011111111100000111100011011101111101100110110100010001100100010101011000001101000010111110011011000100100101010110001011100101110101111010100000110010011100010110101100110100110101101100000000001001110111001101111110000110010000101010010001000110011111110001111100111011000011100110101110011011101110001011100100100001000110000101101101000000011010111011010010001010110000011111010000000011101111010011110001100010010110010000101001110011001100100010110000010011000000101001011101000101101001110011100000101101011000101000100100110101000100110101000101001110100100110110011010111011101101100011100000111111010101001100111001111011111010001011110000010101001110100001111101110010010000010111011101110000011000010001010000110110010111001010001010000011011001101100010100111011001010011010000100100110100000011000000010010101001100011101010001100110000100101010001010001110000101010010001011000100000001110000111001100100000111100011010001101101110100010011111010011000000110001000110010111110011001100001000101011110111110001001111001011011110011000100100110001101010110011000101100011000011111011111001000110100001110110001100100101111011110011011111101010100111110110001001101001010101001100001010000111101001101010100000000000111000111110001011000000001010011000110000000010100001001101110101001010001110110011001000100100000100100111110001011000011100010001110111001111011101010010110111111010010100101011101000101100001101110111110000001110000111101111000110001101101100000100011000111101000101011011100100101110101010110101000110011110100010110100001110011100100100101000111100101001000101110011100010010011101111110010010011100101101111101100010110010011111100001111010010010110111001111101000000001101101111000000110110000000001000100100000011001100111111011110111001111010110100100110100111011001111101011111000001101101111111100011101101001101001001101000001000010000110010100111000000000000101001101010011111010100101001101010001111111100000110111010011100000110100101001011010110110101111011110110010100110010101101001010111111010001000010101000010010100011110100010101010000110101011110100101011001100010000011110111010001111110000101001101111111010000111010000011011101001101010111101101011111001110011010011011011111010000000010010100101101010 : 0)))))))))))))));

    parameter SEED0 = ((WIDTH <= 64) && (TYPE == 0)) ? 64'b1110110110000110101010111100101011110101001011111001010100110000 :
                     (((WIDTH <= 64) && (TYPE == 1)) ? 64'b1010101010011111100011011111010010111000010010110100100011010011 :
                     (((WIDTH <= 64) && (TYPE == 2)) ? 64'b1111010000100001110110000001100111110010100100001010100100000010 :
                     (((WIDTH <= 64) && (TYPE == 3)) ? 64'b1100000111001101001011001001100101100101001000001001011101001010 :
                    (((WIDTH <= 128) && (TYPE == 0)) ? 128'b00000100100000011010011111110010001110010011011101001101010011101010101101000101001011001010001000001110101011100001000011111100 :
                    (((WIDTH <= 128) && (TYPE == 1)) ? 128'b11111111010001101001101000011000000101100100000001011011001010011111000000100100100101111010000111011000110100010000101101111110 :
                    (((WIDTH <= 128) && (TYPE == 2)) ? 128'b01101011100010000100000100011111110111011000001001110010011100101101000000011001010010100010100100101000111101101100110010001011 :
                    (((WIDTH <= 128) && (TYPE == 3)) ? 128'b00000010001000010010110100100000111011010001101010101100101100011001011001001010111010010101100101011111110001101011000000101010 :
                   (((WIDTH <= 1024) && (TYPE == 0)) ? 1024'b0110011010101000110000111110000010001010110100001000101000100100011000101101011011000110011100001010101100011010010000011011000101100011011110010101011011000110011010000101110110010001111001111011000001100010010001111101111011010010111001010000110000010110101010110111111001100010001000110011010011100001101010110101010000011011001011111001111010110010100010110101001101001100100000010111110000000111111001100100110010111000010001110111101110111101110110010101000100111011100101100011000100110000010101001010000011100100100101001000010101010110100010100011010010101000110110010010010001111111000110000001110110110010000001011001111111111000011011111000110100111010000000010101101101001001000011010011110101101101101010011010101110010000011001011100001101010001011111100100111110000011001111110110100011100011101101101110101101001101000111111100111111110100110011000011111111100110001101001001000011011100101110101000011000010011010000001110101110100001011011001110001000000000011011010110001001000101011100000011000001111101 :
                   (((WIDTH <= 1024) && (TYPE == 1)) ? 1024'b1010100100000001111111010111101001001111111101110101101010011110101101001110010011111010001000001011011111010011111110001000001111111010111011101011101111111100010100111000101001001110110010110011000010101010111101110000001000011111001011010111011111110111000110100100010111011011010011011100101001011111100010010011000110111100000110110010000011110010001110100111001000010011010011000011010001100101111110000011110100010110111000011100011100010001111000111111111101100101011000000000101011001000010110000100000010010101000011011010100010010001001011110100100010111011011001111101001100100110011010110100110100001110111011110000110101111100111111100000110000101001101100101001000110111000001100110000010111100101111010000000011010111110100001111101100011010111100011000011111000110111100011100111111101101010011111011100000000110010001110011111010000100000000011110001111111100001011000011000101001100110001100001100001010011111011010000111100001100001111100111010110111100100000100111100111111001000111101111001110001000101 :
                   (((WIDTH <= 1024) && (TYPE == 2)) ? 1024'b1111100011010100101010101101101011111000101011100111110110010110100101000100011111111111110101000010101000001100000011110110000111101010100001001000110001000000101000111111001001010100101011101100101101100101100101010010111100111001001101111101011000010100100000000011010111010001100011001110101111100011001011100101000101101001110110011110100011010100111111111001010110100000100010000110011001010011110101011011011110010101100110011111111011011001011000111011100101000101010000100101111000111000110001011110000010111110001101100000110100101010101000101011111010001001001110011101101100101011001110101111011000101101001110001011001100001100000111011101001110111010010001000001000011010111101001101010000011011111110111101011101001111011111000110110100100011101111000101011001101010011101100111010100000110010010001011111001111101100100100111100011011100001001100011101011100110111111011100000011100111011001100110000101000010010111100100101000100010010111100111110001100000100101001100010101111000000100010100001000101001100 :
                   (((WIDTH <= 1024) && (TYPE == 3)) ? 1024'b0000000011011000000111110010110010010000000101110011111101101101111010100100100000101001101010110111110001011110111111001001110001010011011110011101001111010010000001101110000101111110000111111100001011000101001001111000110010011100100110101000011011100101010001000111111110111000100100000000011010011111000010010001001011000100101011010000100110110101101000001010001000101110011010000100010111111010000110101100001010000000010101011110110011001110001011100111010110101000101000001100101101110100100011011101110001001111111001001101010011000110100011101101011000101011001100100001100101100111111000001110111011100101011111001001100001010011011100011101001011100011010010110100100000111110001110110010001011100101110100010001101000111101001011011110001000101010110110110011100100001010100100110110111101011100001110010010011110110100111011000111001010011100001001011111011001011111000010111001001100111110010010011101011010110100000010110010010111001111010100001000011011011111111000100101100010011010111110011010100110010000 :
                   (((WIDTH <= 4096) && (TYPE == 0)) ? 4096'b0010110011011110111100000101101010110000000010010101111101011111011011000001100001101000100111011010010101110101001000101100101000000100101010110010100110100100011000100011101101011110111000010110001000001001110101001111100010010011000001100100111010000010100111001011101010010010001010010000111001010011101000000100110100010010000110101010000010011001001010110111101000000011010110001101101101100010011111100101111101011000111000010101000100100100000000000001110111100110001011110001110000100010010101111001010111010010001010011010010111111111001010001011101110011111011001011111010111011100010101101101111010011101011010100100011110110111101001011110100111101000110100101010111011101110000000101010000001011000101101000000010101110110001011111101011001001010011001000101110001110010001001111101001100001101011110110011111011101101111100101000010000011100101111000101001011000001011111001101110111101010111111111101011001111011010010100100011111110001110011110111011101001000111000111101011100100110000111111100000110010110000110111011011000100111101010011111011100000101010100101110000111010011101100001111111110100101010110000001111010100110111110110100001000100100001110010111110100001100001111000100001010000000010000010001111111001110001011001101110101010001001100110000111011100010010110100000111101101001010111110010000001111001101111100000100111010011111100100100000100011110011011111101111010010110001111001111001000000011110000101110111011011011001100011001101110011111011011001001110100100011100010001011101010110001011010100011111011001111110000100000110011001011001010101011011001111001011011001100110101011001101110000110001011100101001100100010010111010010101001101111000110111110110100000000111010100100111011000110100000011011001111100001000111110100101011110101001100001001001100001110101101110110111001100101110110110101010110010000100101101001010011110000000111010100110010110001001011111111101000010100100100101010100010010111001001011001100101110001001100101100110101111101110101011000001110001101111101101000010110011110111010101010111011010110001001011011010100010111000001011101011010111000000101100100000101101110110101001101100010110101000011000011111101110110010110111001000100011111011011001011010000000001001010011111010010100011110010001010101000100001000111100110101000000010011101010111010001000010010000001000111110111001000100010010110010001110000000011101111101110000101000111000101111000000110101110100011100111011100101010000011110101110110111000110000010010010000100111001011010111011011001001011010101111110100100111001001111101000010011111101000111010000001110011101111111001001001001010000111100110110100101111000011000010000101111011000000111001010111000100011101110001010000000000000011101110110010000000000111110011000111001000000000011001010011100101111110101011011000011010000101001110101010001101111010011011010101110010100110101000001010110000100101010110011110001100001101111110101110111100111100110011001000101001101011110000101101011110000010001010101101110111100111101001001000110111000110010110001101110000110100001000110000011111101001010101010001100111100110000001010101111010111110000100010001100011001111110111111001110011101001111001001111101010010101010111010110011100111101110111101000001010111000101100011001110001010110011111110111011111110001100101010001100000011110111001011100111001001110110000100010101110101001000101101000011011110110110000111000000001110100110010111011010110110101001000101101001011110111110010110011110101101100100000010110000111100101111010000000101110000001100110110110011001110010010010001110010011011000101100001101111011000101011001101000101000011100101010110001101111101100111000100011110111111100110100010110110110110100110000001011011000110111111100001001000100001000000100000101100111111110111011011001100011000110010111011111110111001111111001001000010111001010001000000011000100110110101110100001010001011011101110011000101110000001101011111110110001111111011100101010000100000001001111110001100011011111011011011000000000100001111111110110101000011101101100001111010111000111011110110011011000000 :
                   (((WIDTH <= 4096) && (TYPE == 1)) ? 4096'b0110110010110000011010001010111000011110101110001001001111001011001101000000000111000000101101101011011001100010110111110011101111000011011110101110100010110100111100111110110111111111000100011000100011111111111000110111000110001011110011001111110000010000010011011110110101100011011110010011000111111000000100011110100101110110100011011000000000101111011101100001101111011000111101111001101000111111001101010011110010010001111110101011000100010001110101101000000110100011111000011000010011110101011010110001111011101000011111000011110000010110101010011101110100000000011001001110000100100001110100110001100011000011111110101001110000010001110001110111011000100011000101110000001101101110100100100000010011110110100110001011100011000111110110111101111000001001100100010101111110111100010000110010111110010001000000000011101000111010000110100000100010111010111001101111110100011011100111010101101011111001100010000010010111101011110001100100110010010011100110111011110101011111011111011100110000001010110100111011000000001010010001010111001110001000001010111111000101011101010111000111101100001011110101100011100100101001001000000100010111000001011101111101101101100101011001111000110001111110110011101101100000001110010011000010011110100100001011110001010110100010101101011111100111100101101010101110101100100110101011100001110010110011100101010111010000001111100010101100000000110001111011101101001100010010100101101100010100010111101001100100101000010011100101000011110100110000000110001100101001000010101001000100111000011010001101110110100010100011010001101100011111001001000111111000110101110100110100110100001100111110001001001001111011011000111101001111010001011001000101110000000111100010011100111001110010111110011010000001011101110110101110110001111001101001010110010010100111001100000000101110001000110100011111111110101010001001100100100001010110101100110100101100101110100000011111001100110100011111010000111100100101111011011101101011110101100111101100111000000111111010100101000000111111110100001011001100100111011000110100110011010011111000001111001001010000010000101101001000011111110111100010011011111101001001000010010100111001100100000011111110010110000010101110101111110100100100110010010111100110001011011010011010001101100001101101101100101000100111111110001100101101110000001101000100001000110110111000101010001110100110101101011100010011001011111101101001000101001000000100010000100010101111011011000110000011001101111100110010011110110000011000010100010011101101010100111101010011010011110110000101100101011100100010101110111001011111111001011111100000110010001000011101101111111011010100101001010100111010100111101111111011100101111110100101111010001101101100000000010101110001111110001101010101101000011100101111110101010110100111100110110101110011011010110110011110111101001110001101111001110010111111101100010110001110100110000111110000011110010101111000000111000000110000101011011000011010000010011011010010010100000001010100010110000000001011000111111101101000011000100001101010100000110111111110001001010101100111011101000111110111111110111010101010011011001110101000111101110110011000010000111111010101000110110001101111100111000001110100001100101101011001011001110011100101101101011111110010000111100101100101011101111110000110011101011110011100110110111111010111011011011100000001000111011010000110100001000101001010100000011001110011110001111010101111101000001110101111100100100011110010110101011100000101101101001110001110101010110010010010100101100000111011010100000010111101100011100101111100111001101100010011101101100100000010110110101000100000111010101111011010111110011001110100111111111100100001111010111110000001000001010101110100111001010100110100010110101100110011001011011100010001101011001001100000011111110100000111001100001101101111100001010011111101100001011110111111011010111010110011110100111001111110110001100011100000001110001100100011011010001101110001011110010010111011000001100100001111011110111001001001101101100001010100110111001101110101010001001110100111100100110001101010110010010110111111011111110110011010000111111000001001010011 :
                   (((WIDTH <= 4096) && (TYPE == 2)) ? 4096'b1110001001100111000111010010110010111111001010100101001111101001001011010101000010001010010110111101000100111011000110011001101101101111011100110111010101001100110000000111100001110011000010111111001010100000010110100110111111100001110100001111010011111101000101100100011110111100010010100100010100001100001000110101110000110001001111100111100001101110111110011100001010100011100011000100011111101100101010001011000110101011111011110011100101000101001111010010000010110011001001010000111110100101111001011110001111100111000101111110000000101111000000000111010001101110101110101100010101100001100011011001100100101100110010010100011011110010000001000000011101000011101011111100001101011100010010110111000001010111000101010001101110000010011011101100000111101011110111000010000110101101101001011010010010000100111011100110011110000100001001010001001100101010100100010000001010010111101110101010111111100011111000000101001001010011010101011001110100101110001101101011101111001001001000110011110110000010011010110100101000001100011101011100001111110110101111000001011100010111111110110100100001111101000001111011000011110101000110001101110001000010111101110001011110001110010011110100110010111110010010111101000101000101011011010100001011000110100101001011001101011100111001101111100000110110000011011001100001011010110000001101100110100010000110111011010001100110001011010100011001110011101011110111010001101001011111000100111111000000111111000000111111111101011100000100010011010100100011001001101010111100111010110110001010000100000110101000101011011000010100010111110110001101110001110010000111100001010100000001000101110110010011101010111001000001111100100000011000111111110101110010101100111001000100011001011100001000000111010111010101010011011011011100111010000011000101100011110010010011000100000110101101100100100111101101011110101111101010001011010011100010110000101000010001001011011101011001100101101100101001111000001010001000010110001100111101001101111111100110110000101010001001000101000001101101010101111101010110100101000001001101011011010001101101000001101110100110001100111100000010111110101001000101101011101111111111101001001011110011101111010110001101100100100111100010000000111100110000000001101011100010100010010111001101111110000110000111010101111010001100101011010100011111100110101000011101111110110011101001101010001001111100011100001100010101011000100000100100010010100101010100100111111111100111001111010000010110011101110101001001010001110101101101010001101010010000111000011000100110000101110101010011101111111110010000111011110010110001101000011010001011000110100010010111110001010010011110011110111101110101010000100100110001110010001100111111101000011001000010011010000001000011111101010010010011101111000110101111111000011100110011011111010011111000000111101011011010111011110101111110001001101011100010010010010110000100011010011111110100000011101010101110001010100000111101100011110101000100111110111110100001100000010110111000001001110101000011001101010100111000111000010110010010000111111011010001011011011011011100000001100101100010011001100011110111000000011011001111110111001011000011011110011111001110000000111000001010001100011011110000011100100011011010011000010110100100011010111011000111011010101010110101000111101110111011001110010000111011100111100111111011000011100110111111110010011000111011010101001101101011011010000100000011101010110110010010010000101011111100100100001101101101101010011111100000101000101010111110100001011010001100111100010110110011100100011100001111111000110011100111000101100111000001000101101100001000001001101111010001011100000001010001101000100101010100100001100110100110010110110111001111000111010000111011010011001000000001111100011101010101111011101110101100001010101101000010011101101001111010000101101101001011110110101010011000010110111010111101000101101111111000010011011101111000101100100100000011010101100001011111100010001100001110100001110101000100000011101101110001011000010000011011100110110011000111111111111000100001010110111111101011111010110001111010111000101010001010100001110111110010111011001011001011 :
                   (((WIDTH <= 4096) && (TYPE == 3)) ? 4096'b0111000011000010101110101110111110010111011010110111011011000001001000011011100110000000011000111110010100011011111100110001000111001011000111010100001001010100101101110100011110101100111111011101000111000101101010111011110011011011000101000011011111001111111101101000010001000100011110111010000011110000110010101001010011110111100111001001101110001011101111011101110000001110110110011101001011001000000100010100001000101000110101011110101110110000100001011110100110000000011101100111001011001110100100001100010000110011011010110001000101000000011011010011001000111110101001001110110100000000101100000001011000111111101100100101010111010100001000111000000000101010110010111010011010011000001100001001011100010011000101001110110011110101010011110000100001110110010000001101111010001010100101101101111111100011011101000010110000110101100010101111011100101001101100001101010011100101000001010011011111110111011100100110111100011110000010110111111110111001000110111001011001001100001101010101101101110010011100000100010001000100101000101000101101101110101001100010010000011011110111001000001011000011101000011100100000101011110011100100111011101001001101010011100110001011101010111000011001011101101100001000100001100011010000101100000000011101001111110110000010000101111111100101000001110000011011111100010001101011101100101101101011101100000011110010100001101101001110001001100000110110000111001110111100011001101111101000010100000010000100100000010000010100001100000101010100110111100101100011111111100010001110010101001101100011111100011100011101111011011011110101001101111000110001000001000100110110000001000101000010001100001111110101011011011111111101101010101011110110001001001111100011100010000111001011000010101001000111011001111010111101011010011101100010010011110101101000010000100110100110010011110010110001000110110001011100011011000000101101010001100111001001101110111010111111100000011101011011110110001000000100010101001100101110010000000001111001001101100011001010000000110110110111011101000001011001010000110101110000011100101110000000010000000011000101001010010000000000001001011100000000010110101001000111011000011100001001110010110010110010001010001010001011011001010101000001111100111010100100111101100100110010111000101111111110101100010100110000111100111000000111001101001011001011111001011000001000011111101100001011000001111011101111011101010011110010110011001001000100111110110100111101111000100101110101100110110111111111100101101101110000011001001110000111011011110101100100011101100110111101110101000101101011011100111011011110111011110000001110010101011010101111101000100110000000001111100111101010001001000010101111000010011001111011110011100101001010011110000010100100111011001110011101001101110111010001110011011001010010100101110000100101100101111000100111100111000010100000111110011111111011010110100111000100000001000001111100001111001000101111010101011101010010100101010111111010001001000011000101000001101110000011001000011111101100100001010111100011101101011111010100101000110010111010001101101000000110101010000111000010011010110111011010100110110000111000011101001101010100011101001000001000001110101001110110101000000110000101111000101101111110100010100100010101010011100001111010101110101010110011000000100001000111110010010011000010100011011001011001101111000010001000110001001001101010101110010011011110111100110001110100100001111100001110011011110111001000110100111001000100000000000000000000101100101111100101101100000000001010001100101000100000101100000111001011100101101000101110111100011110000001101101000110110000010110001100000111110011100011101010101110101001010001111100011101110111011101101101100111111111010100010010000101101001010001000000101001111101001010100001110111001001011001101000111000010010110001001110111101110111001100110011101000100001001000000111111110100101110101101100011111010000000101010011100011000010011000101100111111100110011110011111110110101011111101001110110100010010100101100101011111110100100100111100001011001101101101101000000011100010100111011010111001000111001001011111011101111111110111100100001111101100100010 : 0)))))))))))))));

    parameter SEED1 = ((WIDTH <= 64) && (TYPE == 0)) ? 64'b0000110110000000110100100010000111110010101101001111000000010000 :
                     (((WIDTH <= 64) && (TYPE == 1)) ? 64'b0111111110010010100110100110010010011110101110000010101110111101 :
                     (((WIDTH <= 64) && (TYPE == 2)) ? 64'b0011100101010111100010001000001011001011011111011101000011000000 :
                     (((WIDTH <= 64) && (TYPE == 3)) ? 64'b1110110011101010110101000000011101100101101000100011100000001011 :
                    (((WIDTH <= 128) && (TYPE == 0)) ? 128'b01100011100001101110101000111001110111110100100011010011010101100100000100001101101110111011000000000101100011001100001110100001 :
                    (((WIDTH <= 128) && (TYPE == 1)) ? 128'b10100011111000101001100010100100110001100001110001100111011010010101101001111010001000100010101111110100111011101100011011011110 :
                    (((WIDTH <= 128) && (TYPE == 2)) ? 128'b11001010011000001000000001111111101111010101100110101111010100101000110010101100000000111110101100101111100001111101010100010011 :
                    (((WIDTH <= 128) && (TYPE == 3)) ? 128'b00011100001001110001000111001011001101110001100001011000111011100010001101010011111110111101111111000111011101111010101111001110 :
                   (((WIDTH <= 1024) && (TYPE == 0)) ? 1024'b1011001111111100111000000101001001110000010101110000111000000101100000110100110010010010010101011011101101010101011001111100100010010100111001010101000101111010001101010101000001111000100110000001001011011010011101011011000111110110011111101110010010101110011110110000111010110100011101111010010111001101000011110000111001000101110001110001011001010000100010001011110110000110000001010010111110001110000010000000011000001000111101101011000010100000101001100100001100000111101110110010111100101110000010000110010110110000001000011111111101111110110010001110110001011001000100100100010000100101010011110000011011001010011011110010011100001001001000100111110011000101001101000010001111100000100010100011001100101100101000101011000110011110010000101001101100010001101110100010110111010001011011100011101101111001001001100011110101110111100100110111010010111000101111001110010001000111110000101001100000100011001001101010110001010001011011011100010011010010000011001001111001011110000011011011000101110011001100000100000000111010 :
                   (((WIDTH <= 1024) && (TYPE == 1)) ? 1024'b1001111000111001001011111010100011101000111111001000111101101110111011000011000010001011100011110100110011011100000001110010010011000100011111101001100000101110001100110001001111110111011001001001000111100001011011101001110011010111100000011101110111001111001101000100010101011000010111000101001111011011011101000011101011010111101111110010100001111101100001001100010110101010111000001011110000001101101010010011011110110001001011111011010100011100101110110001110110111000111010101001010111010111001000111101101001011100111010000001000110001001010010000001101000111100010101100011000100001010010010001001010100011110101101000001001001111111111110110011101100101100111101011100100110000110010000000111001000111111110110000011100100101100111100110000010001011110100100110011101011111101101010100001000000101100110010111100100000101001100101001010011010011010011100100011010100110010110101011101101011100011100101111011110110101111010101111001111100100101100111000101010011010111010100000011000010110101010110101100111110111001 :
                   (((WIDTH <= 1024) && (TYPE == 2)) ? 1024'b1100100110101101110011000111000011001100100111110101010011111101000001010011001010011001000111111100100011111101010000101100011010000111001110100010110101100100100100001110101000100000110010001011001001000101110101000111011111000011101001011000100100011000111001010111010000110110001011110000000101111011111111101001111101000111001011010001111100100001110100000110110001010001110111001110010111100101010000101101000010100000011110000110010011100011001011010010100100110000101101000110011001011001000100010110001111000010010000110000011101111010010010100010100011101001010001110110100011110100010100000010110111111100010010111100011010101010110101100011100011011011001011110001100011011100101101000100000001010101111101010011000000101000110011111001101110101010100001101001010011001011000000011010010000001001100110010110100100000100101110100011000111011101110000000011001000011110001011001100001101010110000100000100110001100111000100111001001110111011010100001010100110100001001100100101100011011010111000010011111110111110 :
                   (((WIDTH <= 1024) && (TYPE == 3)) ? 1024'b1001110011101011000001101000010100000001111001011111010111110001101011100110100101111110010001101111100111110100010101010000110100001001000010101011110001101110010011110100101001011101001011010101101011000110100101101110110010011110001010011001010101101011000010001110010100111010110011101011101010110001011101110111001010000110110001001000000101101000010011111010110101010111110100110110111100111110111000010100011000001111010101000011010110100001001010001010001001111100011101101000000001111101101111101101100101101001011110101000000010100110110110100000000010010011001001110000001011010111100101001110111101011111100100000100011000000010101100101001001011100110001111100101111000100110111000100100100101110000111001010101000011110010111100000100001100000111000110101010111100010101001001010010101011000101000001100000001001000100110101111101100001010101000111010100011000001001010000000001111000110100111101001000001111011100000000011100001000100110101001110111101010000001011110001111100101000010011010000010111111101111 :
                   (((WIDTH <= 4096) && (TYPE == 0)) ? 4096'b0011110110111101110110010000101011110101111011111010010010110011011111011100100100011011100010001101100101000010111101111110001001100000010000101101000111001011000010111101011111101101110011110000000110111000111010001101111000010110100010000110010110111101010101010011101011110000011001110110010000100011101000001010010100110011011001000100101001100010100001000100011011001001001001010101111000100000010011101100110110001011001001000000001101010100101100110111110011110101000100011110001101111011011001000111111100110010010010010010011001111101011011010000010111110111000100110100110010110110000111011100100110100111111010010111010111111010000100101111000101010100100001001001101111100100000010010101100001001011100110010101110001111110010011100101010000010100100101100000000001110010111000001101001011010010000101111000001101101010000101001011010000001110110000100111101100000000001110111010111011111100000110010001111010000111110010011000110110100110000111110101100111100100000011100110110100011000110011010110100100010111001001000100001110011001110001011101100001111101100110001001001011111011101000101101011011100110100011010000101010100011010101101100110110011000000110101111110000101010111100000001001011100100110100010000001011010110100000100110000011001100001110010011111110101001011101101010000011001011100000111100000010011110101000000110001111001010001000011000010101110011100100100001001110110111011011011001111010001000110011001110101101110001111011000000011011110110000000100111100000101001100111000110100110000011010001100010100010000010000110010011001111001110111011111100100101001110010110100110011111001001001000001110001010111110011111011110000100100110111110000011001001110110101111000000101110110111110001101111110011111001001010011011100100011001110111100100010000001011000010000000011111010010101110110101010001111000110010011100111011111101010111100110110001100111101111100010111010111100100001000111010011011110011110000010110110001011001111100010010000011111100111111100100101100110001011101011001110110001000101101101000100000111101100000110000011001101010111110000101011101000000111001011110011110011101000110000110000110011000001100110100111110011001001000111001011001000101011011001011011001110011111000010001001000011011011010101010010110100110001100000100100011110110000100110100110110001100001100011001110000000111010101110010111011001010001100111011100001010110111000110111101100111111111111100100010100110011011110100101010101101111101000111100110000100000000011111000010011000000001001011011010110101100101100010000000111011111001011000100001001100101111000100110001000010111100011110001110111001001111010111100100100111011101001110110001000100100101001001011010001010000111101111111101010100100001001110000000010010000110000101101100001110101100000100000110101011011111101001010100011000011110011001000110110010011110111010011100010000001101001110100010000000100001100001010111110011101010101011110000000100111000101111010010001100101010111001011100110000111101010000100100000000111001011100000010001110111010011101010100100101100011110000111010001110100111011011110010111011010101010101010001001110001011110000100111100001011101011111010000111011000111101000111101010101001000100100100111001000100100110100011100100100111011000101111111111111100010011000000011000101110101011011010010100000010111000101100000101111100000101011110111010100110001100100101011111010111001111111000000111100100101011001000110001110101000101101000010001011111011001101000000001101110001010011111001000001001011010001101100001111100111001000111000001000101110101010100011101010011111111110010011111111010001001000000010010110110110010100001010011011101000001010111011111101111010011001110110000000011110110101101110101100011111011110011111110010011010000100111100010010011001101100010010110110010101110010011111010000101010100100110001011001101111001111101011110010000010011110010010110000011010011001111100110000101010000000011010010111110111110010010110000101011011001100001101000101111111101101011111001101101110110110011000100011000011001100100101101100010011000000110010011101 :
                   (((WIDTH <= 4096) && (TYPE == 1)) ? 4096'b0000101011100101000010100000001001101100001100100010111011011011001011001011111010100011100011011111111001100101100111100101111010011010011001010001011110100001000010111100111001000100111111010011001101001001110010011001010001100001000111100101011111000110110101110110011000110001100110000001111011010101100011011110100100100110111110111000111000101001110011000111001110111111110101011100100011001001111111000000111111000011011000100010101001011111111001010110010100100101000011011001001111110111011100000111011101111000111001110001110101010011001011011001011000000101110001010111111101000100100000011101000000000000010100010010101011011100010110010110011010100101011111010011110011000011000000000100101100100001100001111010000101000000101011000110000011000110111001000111010110010000110000010011000100001001001010000100001101110110101111110011011010101110001011111100011111010111100001000010011110110101101000100010110011110110101101000001000011111010111010100010101111000110101110100111100111110110010101111110001001011110010110010000100100111110001010011011101000011111101010110000110000110101100101001010100001010001000100011001111100010100111001010100010100101101110110110000000111010001011010111101110111001110100110100101001101010100000011101100010101100100110111101111001101101110110000001010011110111010010010001110010001101110111100111000111010011110110011010010101001100100000111001001010010000110110101110111100000111000100001110011110010111101101110000101101000100111011110110110001010100111101010101101001001000001000010111100101000010101010110111011100101101010011100011101001011011101101101101111110010100100011000011111100010100010100001011000000000110101110110111111010111111111011111010010111010011011011000100011001011111011010011101100001010010001001000001111000011111000111000011111011001010110000111010001001001001110111100000011110110011101101000110001011000110100100111010110010011111010101101101010011110111001011111101001100001110011110111110010101110000000011011100010000100000111010001110111010100110010101101101111110111100000010010101111111110110110001110010011101101011011111000001001011001110011111000100000001110111011010000101011101111000110100110010110101100010110111011110001011010000101001000101010110110001110000001111010010100000000100111110100100010011110110000000010100011001110111100100110000000010001010011110001010111011110100001110111100110110010000000010101111100000010011110011010100011011110011110100111011111100110010110010011010010111111000101100100100111001100001101011000100100110101011001110001111110000001011111100011011010011111101001101101010111101100010101011001101101000100110101011101010101011110001110001110010001111110000000010101001110001010100001010101010001001001110000001011100001110010000001011000000001110000001011101100110000111110100011000000111100011001100111111011001101111011100101000000000010010001000101000100110110010100101110000001111000101001010101111101010100111100100110010101100111001101011011111010000001100100010110000111110111110001010110000000111100010110101001000001010111010101110110010110000111010001011001110001101101011001100011000110011011101001110110010001100100001000101110110010110010111010001010100110001010010100011000011101100111010100001011101110011100001111100110010110101011100011111010001110010010111010000101010111011111100110000111101111101000111100110101111110011011111001110100101010001011001000100001000001101001011011100100011111101101000010111111001010100011010000111000010100010000100111011011101001000100101111001110110000000110000101110000101100101111111100000010100001110101010101011111011110011111011111101001111100101010100111000110110001011011011010011110000001010100111111011011011001111100011011100000001000000001100001011001111011011011000111110110010011110010011010001111111100110101110001001101110101000000100001100011010110110001101101111011011000101100011110001111111110000100011011001110110110011011011100100100111001010100111100101001100001001101000010101000011001110111011010000100010101010100000000110010011100001001011000001000110011011110100111110110010010101001100000 :
                   (((WIDTH <= 4096) && (TYPE == 2)) ? 4096'b0100010101010000110111100101011011010101101000101011111001000010100001010010011110010110111100101101001111010100010011111011010111100010111000010111110111110111000101010100001010010000100000111010001101000001101000010010001000111001110010110101001111111011011100011110110011000010001010100001000010011011100101101110101101110100100011100011000000000101101111100000000101011011010101111111111111011100100101110101000000100100011010010101100000001111111010000010010001011001011111111010111010110010111001101011011001101101100011001111001001001111011111100010000011101111010110011010001010011010000111000101101111001111111110000111000110111001100100000110000000011101000101101110000111100111110010111101111010001000111100111000010101100111000100010000100001010111110100000000010111011110011010001000110111100010111001100011100000110011111000100101011010110010101001101111010001000111100101010100100111011011100101100101100110110110011111101111000000111111011000011011111011000010111011100010001101110010100111110000110001010001000110101110111001101101100010011000100111011110100000110000110000101001001110011101111001110001111001111011110011100111010110000010000010001001101100100110001100110101001110011100010001111000001010001110011111110110001110011100010100110011101000110000100001000101010111001111100101100111010111111110011111001000011001110010000000101011100001110111000001111101000001110000101000110010101011110110111110110001101101001111111001100001000010110011011110100110100011000110110101000001001001010110011010010011001001010011010000101110100000101110000010001110011100011010100111011110110011011111100001100111110111001111010100111111001000000100101101101011010010101010000001101001110110011111101101110000111111100011111011011010001001010011000001110010110001010000111000001111000111110001100110000011101111100111110110111010000010100000011000100100001101111010110001110101111110100011001010000000101011001000010011101100101100100000010011000000011111101000001010101111111100011100011110010000111110010100110011100000001001101111000100100110110000110001111011010110000001100000101000001111100001000001101100001101111101010100001101110010111010111100011111100111110101110010010111011110111100111011000101110010101001010000100101100110111110110001011111101111001000100010101011011001100011101100001111110101010001100110010001011101100010110110101101101011010011100111000000000111000111111100011101001010100110000010111001000100110100101010001110100010110001101111101001101000010001011001001011011101101011101110100100101100100000001110110010000000100111110100001001001010101100111001111010111101001111101011000100110110000000011000010010100011000101010111100111000101100110101111010010110000111101011111000100101001011011110000100110110000111011100101011010100000110100010110100101000010101010001011011011001011110101000000111100110011010110101011011111110001001010111110001111000101000101111010110101001100111110100001100010111001010110011000110111101000010100000000110001010110111101101010101101100100000101000001111110111001010010001110111110100111000110011100011000101111000001110000100110011100100110010111111101110111101111011111011100101101001111110001010110101010100100101011000001011111000101111100011010111111001110000100000000011110000111011110001011011111011111000011111010001101100010011111010111111011001110111010110011011111000011000011100010010110101111110001011101101010100111101100000110100000101111110010000110000010101010011101011101111100110110010010110100100010110000011000110001110001100000100001011101001101000000001100001101010010110000110110001010100100100001001101100010011010110101000110101001101110111011011000000100110111011110111001110101000101100010110100011101000011010110111010111111010111000011000010100100001010010100110101010000001011011000000110110001111011101100001111010000001001101110100101100110011101000110100111001000010100000011111101000111011001010110011111110101111000110110100110111111100101001011000110111000001011000010111111000100100101110111010001110000101110110110101001111110111101011100001001001111111011111001011111001101110100 :
                   (((WIDTH <= 4096) && (TYPE == 3)) ? 4096'b1011000100011111110000100011001110010010011101011101110000111010011111000101111010011111100000011000100110001100111101011110000100001111011000101010011011011010110101010101011011010111101001111101110110011000001110011110101110110100111010110111111001000110101010101001101011100000110111010111000110111001000110110001011001001011100100001011001000100011101001111001010011000110010101111101001010100011101110000100011010010011011100110000001101001110011000101100000111100111011000111110110100101110101100100010001111111011000010011000000010101110010110001000111111011000010101000010001111110110111011111010110001100110101001100111000001001001010100000110011000110010101001111000010101001110010110011001001000110000011110010100110110001110100100010010000100011011001011010101010110111110100011001100111101100110010111001111010101111011110000100000101110110001001100001010101000101011011000000011001111011111010010011101100111100111100101110101111001111100101100101001110110110011000001011111010100110110101101000100111111010110111110110101011001111100111111011000100111100111001011111100001100011011001011100101000110000101101000000010100010100010010101001110001100100101011111111001000101000111100110011100010101001110010111110010101100000111000000101010100100011111001000011100110100110010010101010011000001101101101110100101011001001011011011001111011000000111010011000100101001000001011011110100001110111111000101000000111011110001100111111100101101000011101010100111010110110011111101000010010101010100000100001100000011101011000001000101001011001101011001110011010010000010000111000000111111000010111010000100010111101001010001101010010100111010100001101001110110101111001011001011001001101101000101011111111111101101100111110110110000111011100100001011101001001011010000011010110110010111011110011101100000011101100110111010111010010001111001000110101011000010111011011111001011110101010001100011101011100010111001101001111000101111100000111101001011111101110111110101100010010000011101101001000010000100100100011110100101111001011011001111101100111001010110001001101011110010101100111110000100101010111110000000000101011111111011000100000000001100001101000110111110001010100000111010111110100000101010001000110100101011001000100100110100100010011111111011011011101100111101110110100111101010010011000100111001011000110011111111100111011100100110010000001111000100100010001110011110110100100000010010111101111100011110111001110001110100000001000110111100010100100111110010101011101000110000110000010110011110000001010001101001100000111000000000101010010101111100000100010111111111011000010011100001110100100001000110110100010101110001000011011011010110001110111101000101100000110110101001011011101011101010011100110100110110011011110000010111001011001110001101001111101100000101101101011111010101100111000100101011001001110110000101101001000000010000110010110110001000000000100111101001000110011101011100111111010000101011100000001100100110110100011011100111010110001100100000000100001010111110010101101000111010010100011011001000100011101010101010000111110000011100010000011011100000011011001111110101001000001111010100001111101011001101010111001110101011011100000111010111000111011110000011111011100000111111000011011011010100110001110011000010011000110100011000110111010000100101100010100110000111010100101111111000111001111101000000101001100111111000000101111111010100000000100111001100000010100100100001000001001111001101010110101110101000110101111111010000000000100111001001001001110011101000100101110001110110011111011010011110111111100001100100100111100001100111001100010010101000101000101110100100111100000001100100111110000100011011010000110000110110111101011010110001101011100110111100111100111110101011101100100111010011011110110100101001000001000101111011100001101100011101111001001011011100010100101110001111101000111010111001000111010101100110010111111101000111001110010001100010111011011000011100110111011001000011100101101110100111000001001100101100110011110100010010001110111010011101001000010100111001100000010111011010100000000100111011101110100001101001101001101010101000 : 0)))))))))))))));

    parameter SEED2 = ((WIDTH <= 64) && (TYPE == 0)) ? 64'b1000001110011101010100111010001001000110001000110000010010001100 :
                     (((WIDTH <= 64) && (TYPE == 1)) ? 64'b0010001011100111000100000101101011110001100101111110101000000001 :
                     (((WIDTH <= 64) && (TYPE == 2)) ? 64'b1001011100110000101011100010000100111011000111101000101011001010 :
                     (((WIDTH <= 64) && (TYPE == 3)) ? 64'b1101000011010000110001110011100111101011010101111000111101100001 :
                    (((WIDTH <= 128) && (TYPE == 0)) ? 128'b01000010011010011010001010011111001000000010111111010111110111010100110011000000100110111011010010000101100011101011101011001101 :
                    (((WIDTH <= 128) && (TYPE == 1)) ? 128'b11110110100101000111001000001000111010110100000110000101100001000000011001100111001000010001000000010100101001111110000100101010 :
                    (((WIDTH <= 128) && (TYPE == 2)) ? 128'b10101110101010000001011111101100001101011111010101111110000101101110010000101101001111000010100111000110000111100110000111101001 :
                    (((WIDTH <= 128) && (TYPE == 3)) ? 128'b10000110001010001111001010111110110010100011110000110011011111110011010010101010110010011111011001101111101000000000101110100101 :
                   (((WIDTH <= 1024) && (TYPE == 0)) ? 1024'b0011000111000100011001010111000000101010110110000001101001010001010011010101100011101010111101001111111100000001110101011110000100000010100101010010001011101100110010010011110110111011010111110000010111101001110110010000101000110110100111001101111111011010110001100110111000010111111110111011100000000100100001101101011000111101100111010100110110011100101110010111100000100110101001010100110111000100001001110110000000010011100111100111101010111010111111010110010011101010001100101100001110111110100000001011101001101111101111101001010000010011110110000111100110011110000001001100101111010110100001010101110110010010000010011110110111001000101010110001110111001111111000100110000001111000111011110000011011101011000010110001000101110100000010000010001001101100111111111101110000000001001101011010110010000000011011000001011110110000110011000100000011110000011001111110111010001111010111101001010010111001000010000101110101110100000000000001110000011111000100001010011000110110000001011111010111110011001111000111010100010001 :
                   (((WIDTH <= 1024) && (TYPE == 1)) ? 1024'b1011110000011001100001011000001110010110001000100011001001100100110010100001010101110001000110110101110101000001111010010000010111000100001011001010001010001000100110110001010111110100111011100000110110100111011000011111010000010100111010011101011010111110101000001101111000011101000001010100100011100111001011100010100000101010111101011110001011101000110011111000101001011010001100010101100011000001000000000000010010100000000000101110010000011011000010100111010101011101000110010010101100000010100110111001100010000011001010010101010111000110100110010110100000001000100011110101000100000100001000100110000011111101011011010011001011110100010110111101110110011001011000001010111001101000110110010010101100100010100110000000100100111101101000100110110110101111110101110000111110110101011101001110011010011110110101111010101100100010101010110011111000010011111110000110000101111001001111000110001110100000010001010110010001100110010101111010110111100110010110110011001001000111101111011011100001000101011011011101100001011111 :
                   (((WIDTH <= 1024) && (TYPE == 2)) ? 1024'b0010101010111100101000000001010100010001010110101001101110011011001101111100011101001101001101110000100110101110001001100011110010110000000111000111010010101011001101001000101011110010110010011100000101011101000100101111001001000010001001100011000111011000101000011100000111110110011101001001100100101101110110100100000101100011100010111000011110000010010001001000101001001110100101110101110101100110000000000010101101111100011011110011100101011100110000011101111110011101110100111110111000000111111001110000000110110001111100010110010110101000101110111101011110000110001111101010110110001010101111101010110001000110101001101001010000101110111001001011100110011001110100010001001000101111010111011101011001000001111100010000110000000100111011010100110100111010110100101010000111010010101001110110101001000111010011100011010100101011111111000001111011010011111110011100010101011010111000101100011100100110101110100101111111011101000101011100111111010111010001100111100110001001111010101111111011110111010110111110010000010111 :
                   (((WIDTH <= 1024) && (TYPE == 3)) ? 1024'b0101011110110011001111110100000100110101111111110101010000100010001001110100011110011010101110000010100001111101110101110011100111011100111001100011001111011110100001011000100000011100000101010101000010010010000100101010101100010101011100000100000101001110011010111011111010001000001110001101111001111011000111011101011001101101110110000010110110100010100111001111111011000000100101110111010110001011000111100111010101110101100101010101000110011110111010011111100110101000101011110000110101010010001001011000000111100001111110011010101111011000010010001010100001000101111101100000110101010010010111001001110000100110001111101010110001000100011100100001011001011100010011110010010110101000000010010100101001111111101101111010101101110110010000111001100101000110001000001101001100011001101011000100000001101100011001001111110111110000010111010000011101010110001101110011000100110011100000101110101011101010000001100100011110001011101010010101101010101011001111001101101101101101100011000010000111000101100111111001000110101101 :
                   (((WIDTH <= 4096) && (TYPE == 0)) ? 4096'b0001101101011100100010010111001000001111001111001101111010011010101001001000001010001110100010110001000000101010110100000100010111001001000111110000001000101110100111101111101110011111011110010010010001100010101110011011011010000010101100111111110100101100001100011011001000001111011111011010110000000011111010011101001100111000101001000001011001000110111011010001000000011011101111010010101001001111110100100111101011111110111110101101001101101100001101010011101001100001111000010010100110010111100110000001001111100010000100110101010010111000011101110011100100111001011010110010000111001001110101101000011001010011111111001011111110100110001010110111001010010011110110100001000110010110000000010110011110000011111101111010111010101010100110010110000100100111001011111011000001110110001101101100001010100101100000001100111011011000100000010110010100111000001101101010001110101100101101001010100011010110011000100001100000011101111000000101100100110010000010010110100010011001001110110011011010010011101011000010100111101000000001010010000001001101111010110110011110010101100010011101000001110001110010100100101111011010100110101111010000001011110000101101011010000110000110010110001010011010001000111111011011101010001001011100001111001001101001010011000111010001001100010101001101011011111101111111100111101011100100001011010100011100111100011110011001000001011101100110010000011010101110100001000001001100110010011111111111001100001101101110010110001000110111110011000111101110110101011100001110001101111100000110100010010101101111101010100111010100000101011100111001100001100101001011110111000010011001110000100100000000000100101001111000000010111100000010000000111010000100010001000101001100110011001111011010000111010000010100001010010001001110101010010011011000111100001100110100010010111010010010001110001011100011100010101110011000101110001110110101000101101001100010111111001100101000000100010010110101010001000001101010101100010111000011010000000100010011110110101001110000010110110011010110110010101000111010101111010001111101110010100011101001010110000001000101010111100011110000001110011010110100101100010010001011011100110111011010000010110011001010011001010111110100100011011011111111100010100000001001111011011000010111010111100111101001100000001101100001010100000010101110001111111000111000000101100100010100101111010111010100111110000110110000000000000110111110000010010011110000111011010010001111010111000011110011110010110010000011101100011010010110111100100111110001011101101110001001011011000100011000001010011001011001000001010111001111111000101110110110010001000100011001100011010001000101111011010100010000001110011000011000000110000010011000100001001001101100011010001100111001001011001000111101110111101000111110111010011111111010011010101010111011101111011000001010000011000100100101110101000100011001000111000100110011000101101000100100101001101100010010000100001000101101001011100101111111010101100100001010110111000100111110111011101110000101011001100011100110010100010000001011000100100011011010001101111010000000101100111111111101100100100100110000001011011110000001111111111010111101011110001000111000110011101101010111101010101111010101110111111001010100110101111110001100101101010100110000101011000000111101100001100101001101110011011100110001110011100000010011100101110110011001110101011101111011010001001001100010111000111101110000000100101110110010111011011010001001011001010111001100100011110101101001110111011101001011110001100100001101111110101110100101011010000111110000000111110010111110011111010100010110010000010001101001010100010110100110000000100010011101100000000101011010101010010001100000010001010001000000101010010010010000010000110110110010101001001101001100100100111000011100111001000000011011101001100010110000011101001010100110001111010000010011001011000010111001110010101000111011111010010100101100110000001001110111000100010010110110110011110101111000111100111000010011001001100011000010000101110101110100101010101001111000100101011001000110010101001001001100001001011110100000101110110110000000100100011000110100100001100011010010100100 :
                   (((WIDTH <= 4096) && (TYPE == 1)) ? 4096'b1001101100111101111110011011111101011101001000000101011001100011101001110101101001110111000001111100100010100011001111100011100110000011111110001001010001011010011101111100111011110100000111000010111101011011010010111011000100001010010111000100000000111001011101011111001100001011010011001001010010111110010101101001001011111101100101100010101101010010111000001011010101011101100100001101000001100100010000100010000101001001010101011000101110100101111011110000001001110110000000001001100001100010011111001011111101111010100010000011011000000000111100001001011111001111111110011011010111001001100011110010100011111101010110011001110000000000111101010110000000000110100100111100100010110000101111000001111100111110100110000110111001011000010101111100001010011101010001100001001100001111000010111110110000111101011110000010011101110000110100110101100101011100101111101110010001010100001110111100100010000011111001110111110111010010110001010001110111001110111101010110011001000000000111110001011111101000001111101101010010000010010111011000111101000010111010011110010011101001110101001001011000110100001101000101010010111011011111110100111001111111101000100100100010000010100110100000100100010010000111000100011001100111011101000000101010000110010011100111011011001100110100110110010001010100000100111001100100111010110110111110111101010001100000110001100111011100011100111010000110011101010101000110010000000000110110001001101000010111000100101111100110111010001111000100111001011001111100011101011000101000111010111010110000010101100101001000000110101110010101011111110101000011111101001001110010100110111100010010101111101010101101111001001110111000001011010111111101110101101110001000011001101110101111001100001001000100011110001110001101100010000000110010011101001010011111111100010001110010101011001010011011001111111000110001010101101100111011111110101000000011111110100100101001110010000010001111011100100001101100001011011111111100111101100000011011011110011100100000110000100000001001001010011111011101001000111000110000111101111010101101110110100110001111011111011000010101011011011101010011111001100000011111101101001111010001011000001111011011000111111100110111100101100001010100000101101101000011011011000011010010011011111110110011011011000010100000000000001001001010100101101010111011110010010001110110010010110010100101111010000110010000110001100111100011011101111000011101010101100011010100110100000110001101000010110101000100101101010100100001010000110000110001011101110110001011110100011011010011110000100010110011011101110010001111100010111010001111101010111111100011111100110110000110100001011111100101101001111001000100010101001010111100010001000000010100101101110010001010101001110111000101001111001101110101101110110001000111011101111101010011111111010011011010100100001101000000001101001001001001100110011100111010111111110010110010011011100000111100010100000001100010001001100010011011101101011110110000011101110011011101101001110011100110110011000001100111000001101101010101110001101101110000000110111001000101000001101110101011000000000011010111011000100000110110101110000100101001011111011101110010010001010000110000001000101000011001101000011101111001101100011000000001111011010011101010011010001001110010111000100111111000100001101001101110011000100001000000011010000001100110111011100110100100100001010111010101000100011010101000011110110011111011001011010001011110101001000010011101001011110001111010011101001100001010101011011100001011110010101101111100000111110110110010010001111010101110101000001011000010111001011111110011000101100011000011001110000011000010110010011000010010100101100111111100101110000001011001101000110111111001011100001100101110000100110111001011111010111100111111101111001100100000110001111111000111100111110101011110001111110101000100000011101110011111011111110011010001101101001100110001101010000000110010010000000110010011010110101000111001010000100001010011000110000100110101010100100100011111100011011000001101000000100101110011000010010000100101000011010111011101101111100010100000001100101100001110011011010110011000001101010111001010 :
                   (((WIDTH <= 4096) && (TYPE == 2)) ? 4096'b1011101001000101000110011001010101011011110011010111011001110100011110101010001111001010101100111001010110001011100000001010111110000001100000101010000101010010101101010000010101110101111000010101010000010100000111110010000010100010010110111110100000111010001010000101111010001110110101111111001110111000000101010100011100011011110000010101010101000011111011010101001010001101010001110101000011111111000101101001001101011001101001101101110001001001111010000111100011111010010111101011101111100110100101010100011110010101101001111011000001011000001110000001110011011110100100010101000000001001000011101110111101110010001001111110000000011100010111010111010110011011100110100010110000000001110111100101010110000000111110001111000010100100101000101000111001111011100101000110101010111100101011000111001000111101011100001100101101111111000111010101010101011011011011011100100011111001000000101101011111111111101111110110011001100011111101111111011011110000110001110111000101000010110010110011011101110010101101010011100001101000110110110000011010100100100110010101000001010010000000101111011011001000101011110101101000100111110000101101010000111111110000100110011111101000100111011011000000101111110100000001100110100101001000110011011000100111100111010101100111000010110001010100000101010101010010111101010000100101110100000111011000111001011110010111000011110110100101011110001001000000010110100001011011101100101111101100101110101100010111010010010010010111110000100111111011111011011111000000000011100001000111100001011010111101011100111111011010001010001110011100010010010110110000011001011110101001110010111110111011001101000100011011011100111000010001001011111010001110100001101100101001101001101011101001010011100010010110010100000101100011010111000100001110110011011011010111110000011100010001000000000101011010000001011000100001110010000001101110110100010101000110110011100110000110001100101000010010011111110110110001110000101101101110011110001011011100001100011001000000011110011001001111001101101001001110110010101100111010001010100101101100100001100001110110000101011111011010110010011011110110011011010101101010011110101001110011000101011010010010111011010110001100011101101011001101110110011011010000011011101100101101101100111111100011010000000001000010100011110110000110111000001001010111100000111110100101110111011011101000110000010010111100011000000110101001101000000011111000001101101110011000001011001100010000110001111011011010100100001111011111101010101111010101001100101001101010011011001111111110001110101011010011001011110110010001111001010111110111101000010110000111101010000100001000011010101011110111000100001111010011111111000100110111001000001000001101111100010101010000010000000101111000001111001101111100011010011101111011110101100100110101110111101010000111000001111100010110111100101010011000010110100101011010010111011101101011010011001110110100100001010011100010011110001011100101011001100001011111100110110100001001001010010001101101101100110011000101000110100001110011101111001000010111010000000110101100100001101110000110111000110010111110010111001110011000000111111000101010110001001011111100001100111101010000000001011110001010011000100111010011101100011001011100001011101001010100100000110011011001010000100011011111100011010110010000100000110000010101100001101010101000101101111010110000011110110011011001100101010000010001101011011100000001011100001000101000110100011001100010001000010100110100111010101110001011010011110110001010101101000101011100101000010111000001010001101100110001101110101001111101100100010110101100110010001010001101110111101101111101010011100001000110000010111001110011011000000110111101101011000001111101000010111010000101101100000101011111001000010100110111001001010111111100100100111010110011010001000011101110100111000011100010000011100000000001010101100001111100100011011110110001111001011111010110100101111111101010000011111010100101101111110100000000101010110001111101000100100000101101100011001001000010010011101001000110010010101010001101010001111011100111010100010111100000110100010001110010100110100100011110101111110011 :
                   (((WIDTH <= 4096) && (TYPE == 3)) ? 4096'b0100001100101001001110001101001000001001101100001001100001111101000011101101110101111110011100100100110111011010000110001111010111101011001110010011110111111000101010101000101101110010100110010100110011100011101110011011001100110011110101001110001100100001000101101100000110111100111011100011001111100011100110110100100110111111001011110011001101000101011100011011100111110000111000010001111010101110010010010101011101111101101110001100011010011001101111010011000101100110001001100100000110111000111011111001000010001001011110100110100101000110001101110101001010001100000010110000000000110011011110101101100000000010011001100000011101001000001100011011001100010011001101100101101101000101111111100001010101110111010100001111100001011001101101111110100010010101000000100000001101001000100110000111100100001010111110011010011001100110010101001101001011110011000100110001110100111010010000100000000011110100010000101001010101010101101000111000011100011111101101100000001000011101010000100011001001010011010110110001001000010010011110010010001111010111100000011011001101100100100000111111011111110000001111101111010110010111111000010110011010000011100111111000010011110100000001000000111010001110011101101001001010111000111110011001101010101101101110000010010001000000110101110000110110110100001111010111101010101110001101110110011010100100001111001100010001110000010100101101100110000011101100100111000011010000000111001011001000101111101010100010110111001111011001011110100000100101000011011010000101110100100101100110001101111011000100110111101100010000011010111001100010001100001011011110011001001111111001111010000100111101000011101001100101011011010011110101001000110011101011110010100011000111001110110101011101110011011011000011101110011001111111110011010010000001011101001010010100001100000011001101011001100110011101110111011001010111001000101101100101101110011110011000101011111010001110110101101100011000001100001010101111010111111001001101010101000001011100011100000110000011100110100111010100100111001100100010101110110001010101011101011101001001100110010101111110101000001110110101111100000001100011001110001100000111011011101011010110000110011101101101011110110111100101001100111101001011110101111100110100100100000011000010001010111011101100101011010011100000001010011010100100000101111101010001000011100111000110100011111011010101101001100011000001111101101100110011110110111011011011011011110111100010000011101101111111001000000010101011111110100100001110000100001111011010010001100110100101110010111110100011000001111100010111000110101110001010010000111110011010010000010111000110011100001111001010111111111000011000110100111000100000010100110110101011001110000000111110111010110001100110011110011000100011010100010110011001110100101010000100011100101101010111101001101100011101101011100101011010010011000001000010010101110011100001101100110101001110010011110011011001100001010100001100000001100101100010010001101101011010100000101000010111001101110011010100000110000100001000111110101000001100111110111011100100001011010001101110000111110000001010000100000001101111100100001000100010101001001111101110100000010011101010100000111110101001100110111111101100101011101111110010101100010101111100100010010000011000011001110010100001100101101110000100010001010001010011110101001101110101000000111011111001010111110101001110111111000110010100010010110110101110110000111110011000111011100000110110101101101110000110001010100100011110010000000001000010101100111001000101100111100011100011110000111001100001001001110010110110111111000110001010111111111001111011100011001100110101000100110110110000101100111110101010000010010110110110101001101011001000100100100101011101000110100110101000010001110000110100101110100001110000000100010010011101010001100101010010100100100010111111011111000010010100110001010110010110001010101011010010101011101001111110001001011010001110011101010000001011100111000110110101111101011111010001110010101110110101101010010001011101011010101010111111000010111011101110100000001011011001010010011000000110100011000011110011110001010101000010100110101000011101101000 : 0)))))))))))))));

    parameter SEED3 = ((WIDTH <= 64) && (TYPE == 0)) ? 64'b1001001001001010010011000001110101110011010101100000100010100000 :
                     (((WIDTH <= 64) && (TYPE == 1)) ? 64'b1111011111100000101110001110110000000100000010000010011111000101 :
                     (((WIDTH <= 64) && (TYPE == 2)) ? 64'b1111101011001010100111111111000110010111110110100011101010100110 :
                     (((WIDTH <= 64) && (TYPE == 3)) ? 64'b1010000111101000001100010111100010100101001111110110001101011000 :
                    (((WIDTH <= 128) && (TYPE == 0)) ? 128'b00110010011101110101011001110001101000110110100101010110001111010001010010101100000010101111001001000100000101001111100111100011 :
                    (((WIDTH <= 128) && (TYPE == 1)) ? 128'b11101101000010011001111001010011001100110000010101010001111110100111110101001111001100111110011001010010111101010111011011000001 :
                    (((WIDTH <= 128) && (TYPE == 2)) ? 128'b00011101110100111000000001110101100100100011000101101010111000000010001101101000000100010100111011001011100010011001111010000100 :
                    (((WIDTH <= 128) && (TYPE == 3)) ? 128'b00011111010101001010111010010010010100011110001110110111111110000100101001111000001111010111110111111100011011111011001010100000 :
                   (((WIDTH <= 1024) && (TYPE == 0)) ? 1024'b0000100011011101001111101110000110011000111100010001110100111100000001001100001010110110000011100101111101101100111101010110100111101101101100001000010100101001011000100001011100111110110111000010100100001101110101010100000111011010111011010010110001000010011101011001010101001110111011000110011000110100000001110001010101111110111001100001001000111101101100010000010110101001101011111100001101100111010101101110100100000100000100001000100000011010010000111110101100000110111011000110100101011001111110100000001011010000110110000101000001010010101111011100010010001101010111101010101110001100111101000111110101010011100111111000011110010000101111011010001101111010111011011100000101001110010111101101011000011111000000010100101010001100001111010101000000111110011001010101001011101100100111111101011111100000100111111011111011011001111101001100111001000110001000000010110010111010111011010111110000010111001011100001100011100111001101111011000011101110110011101111111010010000100110110001111000100101000100010111111110111010 :
                   (((WIDTH <= 1024) && (TYPE == 1)) ? 1024'b0111010010101110100010111100101001100000100111111011101011100100100110010010101111000010000001100100010001010011011011011000100110101011011010010101100010110110010011001110100110010100101111011110101011011000110001110100011100100100111110111001000001011000111100110110010101110010010001001000011010001101011001101011110000011001110011011010011100100111101100010110110010010100001001101100011111000011100010100111010001111001010001111100101110101110111111000111001110010011010000010111001010101011100010010011111001101000110011010010101111111100110011101110011111010110110101100011011101001001010111101110100111011110000010000010000110011011100100001000101110011101000001010011011110101100111000111000010110011011000101000111110000011101100100101100001010100101010100000010010110111100110101110011000110111111111100100100110101000100111011000101011111011011000110001001101000001110001110000000001111111101010000111000001010000101111011010111110010010010101011101001100100000101001011111101100011101100100010000000001110101101 :
                   (((WIDTH <= 1024) && (TYPE == 2)) ? 1024'b1101100011100111110000000001100110001111010100101100111000001100000111001101101010111010011000110011100011100110001110000111000100010101101000000011101010101010110011111101011101001011011011010110101000100000101000000101010101110001101101111100110001100000110100111011000111011010010010000111011111000011000110100001010011000001100011100101100111011101100110011101101100010010010001011101001011000010000100111011010011111000111000010111010110010110010100110101111010100100010000101111011001011000101111011111011111100111000111101100001101111111001110000001001000011011010111010001110001100011100101100101100101010100010011110011011111001100111011001100100111111111110101111011010110111100011101111111101111001100101000110100011000100111001101100011010011101100111011011001101001001000000111101110000110101010010011101000010000101110100011101111100100011010001100100000101001101001000010000110100000100110011000101010111100000010001111100110111101110001011111000111111110000111111011000110101100101011001011011111010111111011 :
                   (((WIDTH <= 1024) && (TYPE == 3)) ? 1024'b0100110111111001010100010101100001110110110100110010010110001001111001100100010111001101011111100110011010000101011111011010001111010100110011100111101000101001010111001010100000010000101011100001110110110101010001111010100000011010110110101111110101001000111110101101001010110000001100111110101000001011110010110000011000111111001100010001101001011011001000001011001001101101010101000000001000000010011110110111010110111010001100100111111000111011101110001000001100011000001000010001110111111001100010111010100100101101110110000001000100010111010100101101001111011110100111011011000100111111110100101100010100111100011000101010111100010110001111111010010000110000101111101001110001010110011001011101100011000111111100110111011011110111100001001000001011001101010110011111101111111011101000001101001001110000000010110111110000000110100100101000101011000001000110001101011011101000011101110110101011011000110000011010101101001101110011110011111001100000111001111011001101111100010110100110010111001100100111001100010101001000 :
                   (((WIDTH <= 4096) && (TYPE == 0)) ? 4096'b0111010011100010111110100010110001100011101000000100011010001111100011011110000010001011011010101000011011000111111000001110100110000001111011000010111011100110101000000010001010010011101101100010110100010100100111111001111101010111001101000011000111111100000100100010110001100110011110111001100101100101100000011100011010000010000111001011101001001011101100100100011001000001111101000000101111110011100100011111001110001101101110010100000000110101101010001110100101010011011011000100101000010101111111000010011101010101001011100000101111010000011001010100111001011111101111101101011100000010000101000010000111010010110100000110011100100101001110010100100111110110011111100001101110001001000101100110101001110110010011110010110011001110111101011100111100000100010110010101010010100100011100010001001110011111111110011000011000100101101000001010011111010000010110100011001011100001001001111110111100010110110100111011110010111101001001001010101000101110000101100110101111000001001001000111011000101110101110100110110001000011101000001100001000011010101001001000111100111011010010101110100011101001001110010110110110001100011011101001010001110100010000100100101011111011101010101001101101001100111111111111111100110111000100110010011110001011101000001111000001100111010110111000010111000001010001100100100011011000100001010001111100101000100101101100111001010101100110111011101110001101110000000111100101111110001100001100000101101101111100001001010001011001111110001010100010110110100001011010010111000011010010111000111101010100110111000000101111001011110010011101110000111110001110100000101110100110000011000010001010000001110110101100100101111010110000100110100000101100100101000110011111101110010010001100100110110101001011010000111011010011001100101101100110000011110011100001001010111011001001000001101000101001001101001000011100111001011100001001101011010100100110011010100110011100011000101010000001100001101011101010110011100000111011110110110011111100101101110100010000000111011011100000000010110000011000011001011110111000011111111100101110110111100110110100011011110001001010101011001111001000011001000110100001001100000011111011110011000111000011101100100111000101110001000110110000110100110000111101001001110000110001000001000000101010111000101110101000010001111110101000100100110011100000110001100011111011000100110110011001101101001000010011110100010101001111101011011101000011101000001011001101010001000100011110000111110100110100001000010110010001001000101101101010000100111110010011101001100101111101001110111101010100101011100110110001110000000101001111001011011001111100111111011110100101001000011100010100110001111101101100101110111011110010100000111000000010010010011110000011010100111001001011000110010010000110100101110011000111010010000101001011100000000011111111000011000001101001010110000100011010001011110011010001101010110111001001111101011010001100111011001000010111111110010110010110110100010100111010111000110000000110011011110100001101100111110000000011011011011011111000100101001101101111101100010111110111111011001011000111000001010011001101111111011111001111100110101001000111010001101101110111110000011010010110000110101000111101101001001000011101010010111010001101101111100011010111010001010111111111000101100110001100101011011100000111010011010010101001001101000000000010111110100000000100000001011111000111100000111011000101110000010100111110001111111011101011100111010101001011111111001110000101000011010001110111000100100010000010110001001010111010111010010111111110010010100110100100111111011011110111100111001011000001000101100110101110011101001010010100011000110001000100100010100111011101100101001001100111010000011001101000001010100101111011110110001001101001010110111010110001000100001101110100010011011110100001001100000111101101101001001101010011111010001111010100110100010000010011110110000000111100111101000111111011110010010011010001011000101101111001000100111011001100001100100010110100010100011101100111111010111101010111001011110001011000010111111000111011110111001111011101100011101110001010001111011010001100110001110110000011000010011001 :
                   (((WIDTH <= 4096) && (TYPE == 1)) ? 4096'b0100110000111110101001000101111111100110110111110010100011010000100101101010000000111111110010100111001100101101011000110101001101100101001100111111101011111011011001010101100111100010100101111100110111110000010111111000101000110011111010111011000111110011010000111110111000001001101110111000101100110000010111011001010010001011000100011010011100110000010101101101000001001000010010101011010100000001001101111001100011111100010000110010101000101100101100001011100110101101001001111101011100000101101010101111001011011001111000001011011111101100010010110011111110001011110100100010001110110011110111101101001100111110010100001001111001010010010110100101111110111100101110111000110111101010100111011101110110100100111011110000101101000001100110100110010001001011000111110010001001010100111011011111101100000000111001100111010100111010010110001100101000000011011001001110110000110100111111101110001011101000101111101110010000010100001011001101100001110000110101101001100110101011010101011100100000100111001100011001111010001000110100111011001011011000110001001100110111010101000000000010101000001001001010110101011110110111010111011101000000110100100101000000100110101010011010110100101110100101101111000011010000100001011110110011011010011100010001000111011110111011100001010011100011011101101010000011100100001000011100100001010010101101101100111000001011101110010010100100110010111011000101100111000001011110001010001101110101011011011101011010100111110010101100011001111100111110111111110110001010101101110001101100101101000101110101101000110000000000011101111111001110111111110101011110110010110000111011000011110011010101101101010000000101001110010010111101011111000110110010011101010111000000001011100010001100010000101100100100010101000011101110101111111001011010100111000110000010011011000000110010010011101000101100010111110100111000000000111000001100011000011000110011000101001010010110011010100100010010110010101100010110001011110101101000111001001111100010011000000010111010110110111000100010000001100010110001111100001101111100010101110110100010000001001001000101101101100011011001111101011010001101111011000100100011101100001100110111011110100010110001101100100000000111111010000010010111011110111111110101110111111011101111111001000101010001101101110011111001100001000101101010010001011111010111000010001010010101101011110010110100010011001001010010001111001100011001011010110000011011001111110100001111110101000001100110001011010010110101010101101101110100010001111000011000001001010010100001111100011101011011011010001101110000011010001100110001110111110110001011110101111101000110110000100100000110100100001101001001001011000101101110111000111111000010110110011001011000010101000101001100010110000100111001011111010111001110010011011010101001010000101101111100111000110001001011011111010110000100000101110101001001000110011110100111101101111011111001000111110000101001000001100001011100011111100001101010000101110111101110100010001100000000100111100011111111100100011010000100000111111011100011111110111111000110011010011110101001110101110011101001000001000001011111110011001001110011101000001110011100000111000000010110111110111010111001101010110111111010100110101100101010110010001111110001100000011111110100100100010110101100010110010000111011111000111111000110101001100110011010001110100100111000101101011110110100110000110000111001110000110010100001110100000100010000011110110001100101011011010010010010111001100011101011011010100111111001101101100011101010001100001101000100101110101100110011101000100010111011000101111111001110010011001110001011101011001010100011010101010010111111001111111101101110100010100111100100010101110010011001000100000010011100101010000011100001011110111001110100110001101110011011110110110000001011110011010011011101101000111101110000110011010101010011011100111110000100101111010010000110010111111101111101001000000110110100000011011101111100100111100100011111100101100101110111001001101101101000010000100110110001111111111100101111010101001100100110011011111011001100010110101011010110111011100100110000010100001010110001010001111001110001010000 :
                   (((WIDTH <= 4096) && (TYPE == 2)) ? 4096'b1001110111111000101000011101000110100110111000001000110110000110110111101111000001110111100010111000011101111100001001000110110011110010011000111101110011111010101110110110101000100101110010000110110011000101011100110110011110011110110110101011100001101110010001000100001010101110100100101111101010101111000001100110010110010010011001000011010101001000010111011011111011101100100011110100011010110110111101010001001111010101000101001101101110011101001100011110111001110011010011100000001110000001011110111000000101111111110011110000000100000000100000101101000000001100000000001001000111000100001011010100000001011100100100111111111100000001101000001111111100111000111000111011101001001000010111110010011000110010001100000010010100000001000110100001010111010001000011100111010101110001101011010011111100011111000100100001011101111101110100111000010001100000110001100011100100110101001101000110011100101011100101100100000110100000100011011011010001110111000110101101111101010101110000010100110101110101100101100110101100101011110111011100010110100001010110011101001111011111001011111000001000101100101001111111111001011010010101010001110000111001110001000110101000111110001100000101010111111100111111001111110011011101101011011110011011100111010011101111110111010100011111000110010011011110011000000111100111001010110010011101001110011010011011000101010001000111101110111100011111010000100001010001101000011001000011000001110100000101011001000001000000110000100111101011100110010010010110101101000010110100100000001011110010000011001111000011111111000011000110001111111101001011011000000000100011101010100101001101011110011100100110100110101110001010000100100110111001110011111011101110111110001101001110010011101010100000110010111010011011010101100100110011111110101101000100111001101000101100011001001101000100111001010001011001011100010011100011011100110101000110010100011000001101001101000001111111001011000001011110010001101000100001111000000011010011101110000001110110000110000100110011010010000100010100000101011000011010100100000110001100011101001101010001011011100101100100101001111101101110000111010101000110011101100001000101001111011000111110100011001101001111101111000100001111101011001100101111100111010101100100010000011111100100100101000110011110101010101010000001100001100101100000000110010101101011100100001000011100110111001100001001100011110010000111000111111110011010001001110011010011110111000001101101100101000110010111010001101111101110100001111100110010111000101001011100001010111011101110111110111011111100000000001100110110110001000101110101001000100100100110010101111110010011111110000010110100001001010011111011110001111011001101001001111010100111111000101001110010100010000101111101001111110000011101100100001111001000000011011100101001010110100110010110110111100111111111101110111010001001101000100011000000011101100110100100111011101011011100110100110010101000101000011110100001101101100110001100010110011101111000011001100110100000111010011100001101101110111011100101110011000100110000100100101100101110111111100111011001001100100001011000011101110110110111011000011000011011011011111101001010011100101111100110111100001110110101101100000001101001010010100001000111100101101111000001001111000011110111100101101010000000100100011000100011101011000110110110101110001110111110011010110111001010110001011001001011111100001100111000000110000100010111101010111001101111001111011010110110101100011011110100011011100100000110000001110101000100111010010000101110111111011010111011001001101101001111110101011011110111001011111101010010111000100111100010110000011001011110100000100011011100110010111111001011111110010111001110001001010010001011011000000011100000000111100111011011111001000011000011110011011100101110000101100001000001010100010101001101100100000111001100100101110001000000110000111011000110001111001100000110100101110110110000000010000101110001111001100110111000011101010000101001111101011010100010000011101010111011011111100001001110000001010100000101011101100000101011100000100011001110010011101011010000000110011011101001011010110110010100101010101110011100 :
                   (((WIDTH <= 4096) && (TYPE == 3)) ? 4096'b0000001010110101011011110000001000011000000111111010111011111110100110101010101101001001010101101011011000100000101011110100000100011011111011110110110001100000110110110100011000110100100100100100010011110001100001100011101101111010110010000000010011000111101110001110001001101100010000000010101101001101111011000010001010110111110010100011011010111100010111001101110001001011001000001110110010010100101101001101100011111011010100111110101001011111000101011000110011010111111111001101110010001000101101111000011111000001111100010110101111110000001001101100001101101011101011011111011001011100011011011100010111111000011001111101111000101001010001000011110000000101100111111000100011111001111001100100101000001100101110110000001011101101100011100101111111101110001001000111000000101110100001111111110011111101111100001111000101100011111101010101110000001111111111000001101000000010010111111101000110101110010111010011010101010110101001110010111001010000110101000101110110000001001001001111011110010001111110001101011000111000111001000001101101111101001101001001001010000000110111001011000001110000111110110100111010100010110001010101000010100010100001110111010001000101001001001111111011110010111110111011010001101010110100001100111011100010110110010010011001110110101011001001100101000011101101011001110111100111000010110101101110110111111000111000100101110001111100001011110000100110100100101110101011111111101110000001111111101010000001011111000101110000110010110111011110000010001101100000100011110100111101000001001100101010101000001111101010101111010100100111000000111011101110100100010001101101101100101010010001011101000111100011110010011111110101001010100100101000110111110110111100100011110111110011111001010110100011001011100011111011101111010000110111010010101101111000001101000001011000110111000001011010001111111100111010111011000010000110110001101010111011100100110110110011010000100111001101010110000110011001111110110100010010100011001101011111010001000101010111001110110011110110010111111101000001000010010010001000010101001111000001011001110000111001100111000011100001111010001101101010110100011000101111010110010000001100110001100111001100010111111000010111111111011010101011111011010010101000010000110011011100001101011111110100011001111110011001001111110101000111100111111000110100001001101000110111010011111111111100011000110010000000000001001111101000000011100101010101001111100101100100100100101010111001011101100110100101001110001100100101101010010111011001110001000010111100110100110001010111101010111110101100001010011111010100101001011100111111111001101100011110010001010101110000100010100110000000010100100011001000010001011000010101111100111101011001111100101101110110111100110001100111110110111011010011010110011010110001000000100001101001001000100010010000110000001111011011011000010010001011010101011011111100010000000001110000000011110101001111010111111111101001101001000011011110101100110110010010000100000000011000110101001001110100000110011110010001111010110000100100110110101110011101011100111000001011111001111010100101000011011010001111110011101000010111111101110010010110011110010100000101001001010000100011001011110101000101011011110101100111110010100100000001001111110001010011100111100100101100010000010111010111010101010100000001110111110011101111100000010000110011010111011100010101010010101111000111101100001011000000110111110110001001010011110010001111011000101100000010100110010100000100111001001101010110110000000111001100001000111101010000000100111001010101011101001100100110001101011101111010000101000000100111001011001010110000111001101011101111011010100011001100011111100010001110101111001100101011110001101010001101100011100000101111011010111000111110101100001101110001010010111010110000111100000101011111101000110010010000011100100110100100011101111100001100010111100101111111100000010101000000110110100001010001010011001010111110101000100011110110011011110010010000111010111110111011101101011010011010000101011000001111111010011011000000111010000000111111011011010001001100001110100100011010111101011001111011010010000111110101100011011010 : 0)))))))))))))));

    reg [REGWIDTH-1:0] x [0:1];
    reg [REGWIDTH-1:0] s [0:1];

    always @(posedge clock) begin : XORSHIFT_PLUS
        if(reset) begin
            prn <= SEED;
            s[0] <= SEED0;
            s[1] <= SEED1;
            x[0] <= SEED2;
            x[1] <= SEED3;
        end else begin
            if(enable) begin
                s[0] <= s[1];
                x[0] <= (s[0] ^ (s[0] << TAP0));
                x[1] <= (((x[0] ^ s[1]) ^ (x[0] >>> TAP1)) ^ (s[1] >>> TAP2));
                s[1] <= x[1];
                prn <= (x[1] + s[1]);
            end
        end
    end

endmodule